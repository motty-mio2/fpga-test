
module KEY_AND_LED ( A, B, F );
input A,B;         // ??????,??KEY1  KEY2??A B?? 
output F;          // ??????,F???LED???
assign F = A & B;  //??F??1 LED?????
                   //??F??0 LED????
endmodule
