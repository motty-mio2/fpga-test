

module ledwater (clk_50M,led_out,f_led_out);
input   clk_50M;       //??????50M
                       //????????50,000,000HZ
output  led_out;       //???????
output  f_led_out;     //???????

reg [24:0] count;  //??????25000000?? ??
reg [24:0] f_count;//??????12500000?? 0.5?

reg  div_clk, f_div_clk;
reg  led_out, f_led_out;



//?????????????
always @ ( posedge clk_50M )
begin
if ( count==25000000 )
 begin     //??????????????50,000,000HZ
           //?????count??????????25,000,000HZ
  div_clk<=~div_clk;  //?????????0.5?????????
                      //????????1Hz??????
   count<=0;          //???????
  end
else
  count<=count+1;     //??????
  led_out<=div_clk;  //??????????????????
                      //?LED????????
end 

//????????0.5????
always @ ( posedge clk_50M )
begin
if ( f_count==12500000 )    //?????count??????????12,500,000HZ
 begin
  f_div_clk<=~f_div_clk;    //?????????0.25?????????
                            //????????0.5???2HZ?
   f_count<=0;
  end
else
  f_count<=f_count+1;      //??????
  f_led_out<=f_div_clk;   //??????????????????
                           //?LED????????
end

endmodule














